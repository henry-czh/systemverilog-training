virtual class default_gen_cbs;
	virtual task set_default_gen(ref generator default_gen);
	endtask
endclass
