class generator;

	mailbox gen2drv;
	event 	drv2gen;

	int num; //num of trans

	transaction trans;

	function new(mailbox gen2drv,event drv2gen);
		this.gen2drv=gen2drv;
		this.drv2gen=drv2gen;
		num = 10;
	endfunction

	virtual task run;
		repeat(num) begin
			trans = new();
			assert(trans.randomize());
			gen2drv.put(trans);
			$display($sformatf("@%0t: generator\t-->gen one pkt ...",$time));
			@drv2gen;
		end
	endtask

endclass
